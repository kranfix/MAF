/* ADC Reader
file:	adcreader.vhd
author: Frank Andre Moreno vera
e-mail: frankmoreno1993@gmail.com
*/
library ieee;
use ieee.std_logic_1164.all;
use work.mafpack.all;

entity adc128s022 is
port(
  EN_N,clk: in std_logic;
  ADC_SDAT: in std_logic;
  ADC_ADDR: in std_logic_vector(2 downto 0);
  ADC_CS_N: buffer std_logic;
  ADC_SADDR, ADC_SCLK: out std_logic;
  ADC_DATA: out std_logic_vector(11 downto 0)
  clk_out:	out std_logic;
);
end adc128s022;

architecture reader of adc128s022 is
  signal cycle: integer range 0 to 15:= 0;
begin

-- EN_N to ADC_CS_N and clk to clk_out
process(EN_N,ADC_SCLK)
	i: integer range 0 to 15
begin
  if(EN_N = '1') then
    ADC_CS_N = '1';
	 clk_out = '0';
  elsif falling_edge(clk) then
    ADC_CS_N = '0';
	 if ()
  end if;
end process;

-- ADC_SDAT to ADC_DATA
process(ADC_CS_N,clk)
begin
	if(ADC_CS_N = '1') then
	  ADC_SADDR <= 'Z';
	  ADC_SCLK <= '1';
	  ADC_DATA <= (others => 'Z');
	  cycle <= 0;
	elsif rising_edge(ADC_SCLK) then
		if (cycle = )
	end if;
end process;

-- ADC_SADDR to ADC_ADDR
process(EN_N,ADC_SCLK)
  variable i: integer range 0 to 15;
begin
  if(ADC_CS_N = '1') then
    ADC_SADDR <= 'Z';
	 ADC_SCLK <= '1';
	 ADC_DATA <= (others => 'Z');
  elsif falling_edge(ADC_SCLK) then

  end if;
end process;

end reader;