/* ADC Reader
file:	adcreader.vhd
author: Frank Andre Moreno vera
e-mail: frankmoreno1993@gmail.com
*/
library ieee;
use ieee.std_logic_1164.all;
use work.mafpack.all;

entity adcreader is
port();
end adcreader;

architecture reader of adcreader is
begin
end reader;